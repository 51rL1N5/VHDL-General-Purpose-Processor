library ieee;
use ieee.std_logic_1164.all;

entity mux4x1_4bits is
	port
	(
		A0      : in std_logic_vector (3 downto 0);
		A1      : in std_logic_vector (3 downto 0);
		A2      : in std_logic_vector (3 downto 0);
		A3      : in std_logic_vector (3 downto 0);
		SW      : in std_logic_vector (1 downto 0);
		output  : out std_logic_vector (3 downto 0)
	);
end mux4x1_4bits;
	
architecture behavior of mux4x1_4bits is

begin

	process(SW)
	begin
		case SW is
			when "00" =>
				output <= A0;
			when "01" =>
				output <= A1;
			when "10" =>
				output <= A2;
			when "11" =>
				output <= A3;
		end case;
	end process;
	
end behavior;